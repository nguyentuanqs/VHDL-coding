library ieee;
use std_
